library verilog;
use verilog.vl_types.all;
entity subtrator_vlg_vec_tst is
end subtrator_vlg_vec_tst;
